`timescale 1ns / 1ps

module WB #(parameter WIDTH=32)( 
    );
    // 5 stage pipeline
    
endmodule