package global_params;
    parameter int INSTR_WIDTH = 32;
    parameter int DATA_WIDTH = 32;
    parameter int INSTR_MEM_DEPTH = 1024;
    parameter int BRANCH_STALL_CYCLES = 2;
endpackage