`timescale 1ns / 1ps

module HZRD_DETECT(
    input ID_EX_MemRead
    output PC_Write
    output IF_ID_Write
    output other
);
    
endmodule

module ID #(parameter WIDTH=32)( 
);
    // 5 stage pipeline
    
endmodule