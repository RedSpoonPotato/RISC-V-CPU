`define INSTR_WIDTH 32
`define DATA_WIDTH 32