`timescale 1ns / 1ps

module MEM #(parameter WIDTH=32)( 
    );
    // 5 stage pipeline
    
endmodule