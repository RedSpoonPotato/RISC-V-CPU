`timescale 1ns / 1ps

module EX #(parameter WIDTH=32)( 
    );
    // 5 stage pipeline
    
endmodule